module Booth #(
    parameter WIDTH = 32,
    parameter N     = WIDTH / 2   // For radix-4, N = WIDTH/2
)(
    input  CLK, RST,
    input  [WIDTH-1:0] x, y,
    output reg [2*WIDTH-1:0] p
);

    // ────────────────────────────────
    // Internal signals
    // ────────────────────────────────
    reg  [2:0] cc [0:N-1];                   // Booth control codes
    reg  signed [WIDTH:0] pp  [0:N-1];       // Partial products (+ sign bit)
    reg  signed [2*WIDTH-1:0] spp [0:N-1];   // Shifted partial products
    reg  signed [WIDTH:0] inv_x;             // Two's complement of x
    wire signed [2*WIDTH-1:0] prod;          // Final product

    integer kk;

    // ────────────────────────────────
    // Booth encoding & partial product generation
    // ────────────────────────────────
    always @(*) begin
        // Two's complement of x (sign-extended)
        inv_x = {~x[WIDTH-1], ~x} + 1;

        // Booth control codes
        cc[0] = {y[1], y[0], 1'b0};
        for (kk = 1; kk < N; kk = kk + 1)
            cc[kk] = {y[2*kk + 1], y[2*kk], y[2*kk - 1]};

        // Partial products
        for (kk = 0; kk < N; kk = kk + 1) begin
            case (cc[kk])
                3'b000, 3'b111: pp[kk] = 0;                      // 0
                3'b001, 3'b010: pp[kk] = {x[WIDTH-1], x};        // +x
                3'b011:         pp[kk] = {x, 1'b0};              // +2x
                3'b100:         pp[kk] = {inv_x[WIDTH-1:0], 1'b0}; // -2x
                3'b101, 3'b110: pp[kk] = inv_x;                  // -x
                default:        pp[kk] = 0;
            endcase

            // Shifted partial product
            spp[kk] = $signed(pp[kk]) <<< (2 * kk);
        end
    end

    // ────────────────────────────────
    // CSA Tree (Reduction of partial products)
    // ────────────────────────────────
    wire [63:0] S0,  C0,  S1,  C1,  S2,  C2,  S3,  C3,  S4,  C4;
    wire [63:0] S5,  C5,  S6,  C6,  S7,  C7;
    wire [63:0] S8,  C8,  S9,  C9;
    wire [63:0] S10, C10, S11, C11;
    wire [63:0] S12, C12;
    wire [63:0] S13, C13;

    // Level 1
    CSA csa1 (.A(spp[0]),  .B(spp[1]),  .C(spp[2]),  .Sum(S0),  .Carry(C0));
    CSA csa2 (.A(spp[3]),  .B(spp[4]),  .C(spp[5]),  .Sum(S1),  .Carry(C1));
    CSA csa3 (.A(spp[6]),  .B(spp[7]),  .C(spp[8]),  .Sum(S2),  .Carry(C2));
    CSA csa4 (.A(spp[9]),  .B(spp[10]), .C(spp[11]), .Sum(S3),  .Carry(C3));
    CSA csa5 (.A(spp[12]), .B(spp[13]), .C(spp[14]), .Sum(S4),  .Carry(C4));

    // Level 2
    CSA csa6 (.A(S0),  .B({C0[62:0],1'b0}), .C(S1),  .Sum(S5),  .Carry(C5));
    CSA csa7 (.A({C1[62:0],1'b0}), .B(S2),  .C({C2[62:0],1'b0}), .Sum(S6), .Carry(C6));
    CSA csa8 (.A(S3),  .B({C3[62:0],1'b0}), .C(S4),  .Sum(S7),  .Carry(C7));

    // Level 3
    CSA csa9  (.A(S5), .B({C5[62:0],1'b0}), .C(S6),  .Sum(S8),  .Carry(C8));
    CSA csa10 (.A({C6[62:0],1'b0}), .B(S7), .C({C7[62:0],1'b0}), .Sum(S9), .Carry(C9));

    // Level 4
    CSA csa11 (.A(S8), .B({C8[62:0],1'b0}), .C(S9),  .Sum(S10), .Carry(C10));
    CSA csa12 (.A({C9[62:0],1'b0}), .B({C4[62:0],1'b0}), .C(spp[15]), .Sum(S11), .Carry(C11));

    // Level 5
    CSA csa13 (.A(S10), .B({C10[62:0],1'b0}), .C(S11), .Sum(S12), .Carry(C12));

    // Level 6
    CSA csa14 (.A(S12), .B({C12[62:0],1'b0}), .C({C11[62:0],1'b0}), .Sum(S13), .Carry(C13));

    // ────────────────────────────────
    // Pipeline registers
    // ────────────────────────────────
    reg signed [63:0] C13_reg, S13_reg;

    always @(posedge CLK) begin
        if (RST) begin
            C13_reg <= 0;
            S13_reg <= 0;
        end else begin
            C13_reg <= C13;
            S13_reg <= S13;
        end
    end

    // ────────────────────────────────
    // Final Adder (CPA)
    // ────────────────────────────────
    //CLA     #(.WIDTH(64)) CPA (.A(S13), .B({C13[62:0],1'b0}), .Cin(1'b0), .S(prod));
    //Knowles               CPA (.A(S13_reg), .B({C13_reg[62:0],1'b0}), .Cin(1'b0), .Sum(prod));
    KSA CPA (.A(S13_reg), .B({C13_reg[62:0],1'b0}), .Cin(1'b0), .Sum(prod));

    // ────────────────────────────────
    // Output register
    // ────────────────────────────────
    always @(posedge CLK) begin
        if (RST)
            p <= 0;
        else
            p <= prod;
    end

endmodule
